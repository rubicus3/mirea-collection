library verilog;
use verilog.vl_types.all;
entity Prac4_vlg_vec_tst is
end Prac4_vlg_vec_tst;
