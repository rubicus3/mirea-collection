library verilog;
use verilog.vl_types.all;
entity Prac3_vlg_vec_tst is
end Prac3_vlg_vec_tst;
