library verilog;
use verilog.vl_types.all;
entity Prac6_vlg_vec_tst is
end Prac6_vlg_vec_tst;
