library verilog;
use verilog.vl_types.all;
entity Prac5_vlg_vec_tst is
end Prac5_vlg_vec_tst;
