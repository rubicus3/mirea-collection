library verilog;
use verilog.vl_types.all;
entity Prac1 is
    port(
        Y               : out    vl_logic;
        b               : in     vl_logic;
        c               : in     vl_logic;
        a               : in     vl_logic;
        d               : in     vl_logic
    );
end Prac1;
