library verilog;
use verilog.vl_types.all;
entity Prac1_vlg_vec_tst is
end Prac1_vlg_vec_tst;
