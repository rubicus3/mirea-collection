library verilog;
use verilog.vl_types.all;
entity Prac3_vlg_sample_tst is
    port(
        a0              : in     vl_logic;
        a1              : in     vl_logic;
        a2              : in     vl_logic;
        x0              : in     vl_logic;
        x1              : in     vl_logic;
        x2              : in     vl_logic;
        x3              : in     vl_logic;
        x4              : in     vl_logic;
        x5              : in     vl_logic;
        x6              : in     vl_logic;
        x7              : in     vl_logic;
        sampler_tx      : out    vl_logic
    );
end Prac3_vlg_sample_tst;
