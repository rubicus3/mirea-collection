library verilog;
use verilog.vl_types.all;
entity Prac2_vlg_vec_tst is
end Prac2_vlg_vec_tst;
